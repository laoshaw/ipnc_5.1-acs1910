nameserver 168.95.192.1
nameserver 61.64.127.2
nameserver 168.95.1.1
